module direct_digital_synthesizer(
  input         clock,
  input         reset,
  input         io_initdone,
  input  [31:0] io_A,
  output [11:0] io_B
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] phase; // @[direct_digital_synthesizer.scala 35:22]
  wire [31:0] _phase_T_1 = phase + io_A; // @[direct_digital_synthesizer.scala 39:18]
  wire [9:0] idx = phase[31:22]; // @[direct_digital_synthesizer.scala 66:18]
  wire [11:0] _GEN_1 = 10'h1 == idx ? $signed(12'sh8) : $signed(12'sh0); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_2 = 10'h2 == idx ? $signed(12'sh10) : $signed(_GEN_1); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_3 = 10'h3 == idx ? $signed(12'sh18) : $signed(_GEN_2); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_4 = 10'h4 == idx ? $signed(12'sh20) : $signed(_GEN_3); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_5 = 10'h5 == idx ? $signed(12'sh28) : $signed(_GEN_4); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_6 = 10'h6 == idx ? $signed(12'sh30) : $signed(_GEN_5); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_7 = 10'h7 == idx ? $signed(12'sh38) : $signed(_GEN_6); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_8 = 10'h8 == idx ? $signed(12'sh40) : $signed(_GEN_7); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_9 = 10'h9 == idx ? $signed(12'sh48) : $signed(_GEN_8); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_10 = 10'ha == idx ? $signed(12'sh50) : $signed(_GEN_9); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_11 = 10'hb == idx ? $signed(12'sh58) : $signed(_GEN_10); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_12 = 10'hc == idx ? $signed(12'sh60) : $signed(_GEN_11); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_13 = 10'hd == idx ? $signed(12'sh68) : $signed(_GEN_12); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_14 = 10'he == idx ? $signed(12'sh70) : $signed(_GEN_13); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_15 = 10'hf == idx ? $signed(12'sh78) : $signed(_GEN_14); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_16 = 10'h10 == idx ? $signed(12'sh80) : $signed(_GEN_15); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_17 = 10'h11 == idx ? $signed(12'sh88) : $signed(_GEN_16); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_18 = 10'h12 == idx ? $signed(12'sh90) : $signed(_GEN_17); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_19 = 10'h13 == idx ? $signed(12'sh98) : $signed(_GEN_18); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_20 = 10'h14 == idx ? $signed(12'sha0) : $signed(_GEN_19); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_21 = 10'h15 == idx ? $signed(12'sha8) : $signed(_GEN_20); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_22 = 10'h16 == idx ? $signed(12'shb0) : $signed(_GEN_21); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_23 = 10'h17 == idx ? $signed(12'shb8) : $signed(_GEN_22); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_24 = 10'h18 == idx ? $signed(12'shc0) : $signed(_GEN_23); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_25 = 10'h19 == idx ? $signed(12'shc8) : $signed(_GEN_24); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_26 = 10'h1a == idx ? $signed(12'shd0) : $signed(_GEN_25); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_27 = 10'h1b == idx ? $signed(12'shd8) : $signed(_GEN_26); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_28 = 10'h1c == idx ? $signed(12'she0) : $signed(_GEN_27); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_29 = 10'h1d == idx ? $signed(12'she8) : $signed(_GEN_28); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_30 = 10'h1e == idx ? $signed(12'shf0) : $signed(_GEN_29); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_31 = 10'h1f == idx ? $signed(12'shf8) : $signed(_GEN_30); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_32 = 10'h20 == idx ? $signed(12'sh100) : $signed(_GEN_31); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_33 = 10'h21 == idx ? $signed(12'sh108) : $signed(_GEN_32); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_34 = 10'h22 == idx ? $signed(12'sh110) : $signed(_GEN_33); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_35 = 10'h23 == idx ? $signed(12'sh118) : $signed(_GEN_34); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_36 = 10'h24 == idx ? $signed(12'sh120) : $signed(_GEN_35); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_37 = 10'h25 == idx ? $signed(12'sh128) : $signed(_GEN_36); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_38 = 10'h26 == idx ? $signed(12'sh130) : $signed(_GEN_37); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_39 = 10'h27 == idx ? $signed(12'sh138) : $signed(_GEN_38); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_40 = 10'h28 == idx ? $signed(12'sh140) : $signed(_GEN_39); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_41 = 10'h29 == idx ? $signed(12'sh148) : $signed(_GEN_40); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_42 = 10'h2a == idx ? $signed(12'sh150) : $signed(_GEN_41); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_43 = 10'h2b == idx ? $signed(12'sh158) : $signed(_GEN_42); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_44 = 10'h2c == idx ? $signed(12'sh160) : $signed(_GEN_43); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_45 = 10'h2d == idx ? $signed(12'sh168) : $signed(_GEN_44); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_46 = 10'h2e == idx ? $signed(12'sh170) : $signed(_GEN_45); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_47 = 10'h2f == idx ? $signed(12'sh178) : $signed(_GEN_46); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_48 = 10'h30 == idx ? $signed(12'sh180) : $signed(_GEN_47); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_49 = 10'h31 == idx ? $signed(12'sh188) : $signed(_GEN_48); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_50 = 10'h32 == idx ? $signed(12'sh190) : $signed(_GEN_49); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_51 = 10'h33 == idx ? $signed(12'sh198) : $signed(_GEN_50); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_52 = 10'h34 == idx ? $signed(12'sh1a0) : $signed(_GEN_51); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_53 = 10'h35 == idx ? $signed(12'sh1a8) : $signed(_GEN_52); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_54 = 10'h36 == idx ? $signed(12'sh1b0) : $signed(_GEN_53); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_55 = 10'h37 == idx ? $signed(12'sh1b8) : $signed(_GEN_54); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_56 = 10'h38 == idx ? $signed(12'sh1c0) : $signed(_GEN_55); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_57 = 10'h39 == idx ? $signed(12'sh1c8) : $signed(_GEN_56); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_58 = 10'h3a == idx ? $signed(12'sh1d0) : $signed(_GEN_57); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_59 = 10'h3b == idx ? $signed(12'sh1d8) : $signed(_GEN_58); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_60 = 10'h3c == idx ? $signed(12'sh1e0) : $signed(_GEN_59); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_61 = 10'h3d == idx ? $signed(12'sh1e8) : $signed(_GEN_60); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_62 = 10'h3e == idx ? $signed(12'sh1f0) : $signed(_GEN_61); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_63 = 10'h3f == idx ? $signed(12'sh1f8) : $signed(_GEN_62); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_64 = 10'h40 == idx ? $signed(12'sh200) : $signed(_GEN_63); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_65 = 10'h41 == idx ? $signed(12'sh208) : $signed(_GEN_64); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_66 = 10'h42 == idx ? $signed(12'sh210) : $signed(_GEN_65); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_67 = 10'h43 == idx ? $signed(12'sh218) : $signed(_GEN_66); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_68 = 10'h44 == idx ? $signed(12'sh220) : $signed(_GEN_67); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_69 = 10'h45 == idx ? $signed(12'sh228) : $signed(_GEN_68); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_70 = 10'h46 == idx ? $signed(12'sh230) : $signed(_GEN_69); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_71 = 10'h47 == idx ? $signed(12'sh238) : $signed(_GEN_70); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_72 = 10'h48 == idx ? $signed(12'sh240) : $signed(_GEN_71); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_73 = 10'h49 == idx ? $signed(12'sh248) : $signed(_GEN_72); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_74 = 10'h4a == idx ? $signed(12'sh250) : $signed(_GEN_73); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_75 = 10'h4b == idx ? $signed(12'sh258) : $signed(_GEN_74); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_76 = 10'h4c == idx ? $signed(12'sh260) : $signed(_GEN_75); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_77 = 10'h4d == idx ? $signed(12'sh268) : $signed(_GEN_76); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_78 = 10'h4e == idx ? $signed(12'sh270) : $signed(_GEN_77); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_79 = 10'h4f == idx ? $signed(12'sh278) : $signed(_GEN_78); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_80 = 10'h50 == idx ? $signed(12'sh280) : $signed(_GEN_79); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_81 = 10'h51 == idx ? $signed(12'sh288) : $signed(_GEN_80); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_82 = 10'h52 == idx ? $signed(12'sh290) : $signed(_GEN_81); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_83 = 10'h53 == idx ? $signed(12'sh298) : $signed(_GEN_82); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_84 = 10'h54 == idx ? $signed(12'sh2a0) : $signed(_GEN_83); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_85 = 10'h55 == idx ? $signed(12'sh2a8) : $signed(_GEN_84); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_86 = 10'h56 == idx ? $signed(12'sh2b0) : $signed(_GEN_85); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_87 = 10'h57 == idx ? $signed(12'sh2b8) : $signed(_GEN_86); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_88 = 10'h58 == idx ? $signed(12'sh2c0) : $signed(_GEN_87); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_89 = 10'h59 == idx ? $signed(12'sh2c8) : $signed(_GEN_88); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_90 = 10'h5a == idx ? $signed(12'sh2d0) : $signed(_GEN_89); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_91 = 10'h5b == idx ? $signed(12'sh2d8) : $signed(_GEN_90); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_92 = 10'h5c == idx ? $signed(12'sh2e0) : $signed(_GEN_91); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_93 = 10'h5d == idx ? $signed(12'sh2e8) : $signed(_GEN_92); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_94 = 10'h5e == idx ? $signed(12'sh2f0) : $signed(_GEN_93); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_95 = 10'h5f == idx ? $signed(12'sh2f8) : $signed(_GEN_94); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_96 = 10'h60 == idx ? $signed(12'sh300) : $signed(_GEN_95); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_97 = 10'h61 == idx ? $signed(12'sh308) : $signed(_GEN_96); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_98 = 10'h62 == idx ? $signed(12'sh310) : $signed(_GEN_97); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_99 = 10'h63 == idx ? $signed(12'sh318) : $signed(_GEN_98); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_100 = 10'h64 == idx ? $signed(12'sh320) : $signed(_GEN_99); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_101 = 10'h65 == idx ? $signed(12'sh328) : $signed(_GEN_100); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_102 = 10'h66 == idx ? $signed(12'sh330) : $signed(_GEN_101); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_103 = 10'h67 == idx ? $signed(12'sh338) : $signed(_GEN_102); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_104 = 10'h68 == idx ? $signed(12'sh340) : $signed(_GEN_103); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_105 = 10'h69 == idx ? $signed(12'sh348) : $signed(_GEN_104); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_106 = 10'h6a == idx ? $signed(12'sh350) : $signed(_GEN_105); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_107 = 10'h6b == idx ? $signed(12'sh358) : $signed(_GEN_106); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_108 = 10'h6c == idx ? $signed(12'sh360) : $signed(_GEN_107); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_109 = 10'h6d == idx ? $signed(12'sh368) : $signed(_GEN_108); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_110 = 10'h6e == idx ? $signed(12'sh370) : $signed(_GEN_109); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_111 = 10'h6f == idx ? $signed(12'sh378) : $signed(_GEN_110); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_112 = 10'h70 == idx ? $signed(12'sh380) : $signed(_GEN_111); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_113 = 10'h71 == idx ? $signed(12'sh388) : $signed(_GEN_112); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_114 = 10'h72 == idx ? $signed(12'sh390) : $signed(_GEN_113); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_115 = 10'h73 == idx ? $signed(12'sh398) : $signed(_GEN_114); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_116 = 10'h74 == idx ? $signed(12'sh3a0) : $signed(_GEN_115); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_117 = 10'h75 == idx ? $signed(12'sh3a8) : $signed(_GEN_116); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_118 = 10'h76 == idx ? $signed(12'sh3b0) : $signed(_GEN_117); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_119 = 10'h77 == idx ? $signed(12'sh3b8) : $signed(_GEN_118); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_120 = 10'h78 == idx ? $signed(12'sh3c0) : $signed(_GEN_119); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_121 = 10'h79 == idx ? $signed(12'sh3c8) : $signed(_GEN_120); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_122 = 10'h7a == idx ? $signed(12'sh3d0) : $signed(_GEN_121); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_123 = 10'h7b == idx ? $signed(12'sh3d8) : $signed(_GEN_122); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_124 = 10'h7c == idx ? $signed(12'sh3e0) : $signed(_GEN_123); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_125 = 10'h7d == idx ? $signed(12'sh3e8) : $signed(_GEN_124); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_126 = 10'h7e == idx ? $signed(12'sh3f0) : $signed(_GEN_125); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_127 = 10'h7f == idx ? $signed(12'sh3f8) : $signed(_GEN_126); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_128 = 10'h80 == idx ? $signed(12'sh3ff) : $signed(_GEN_127); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_129 = 10'h81 == idx ? $signed(12'sh407) : $signed(_GEN_128); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_130 = 10'h82 == idx ? $signed(12'sh40f) : $signed(_GEN_129); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_131 = 10'h83 == idx ? $signed(12'sh417) : $signed(_GEN_130); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_132 = 10'h84 == idx ? $signed(12'sh41f) : $signed(_GEN_131); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_133 = 10'h85 == idx ? $signed(12'sh427) : $signed(_GEN_132); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_134 = 10'h86 == idx ? $signed(12'sh42f) : $signed(_GEN_133); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_135 = 10'h87 == idx ? $signed(12'sh437) : $signed(_GEN_134); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_136 = 10'h88 == idx ? $signed(12'sh43f) : $signed(_GEN_135); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_137 = 10'h89 == idx ? $signed(12'sh447) : $signed(_GEN_136); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_138 = 10'h8a == idx ? $signed(12'sh44f) : $signed(_GEN_137); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_139 = 10'h8b == idx ? $signed(12'sh457) : $signed(_GEN_138); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_140 = 10'h8c == idx ? $signed(12'sh45f) : $signed(_GEN_139); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_141 = 10'h8d == idx ? $signed(12'sh467) : $signed(_GEN_140); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_142 = 10'h8e == idx ? $signed(12'sh46f) : $signed(_GEN_141); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_143 = 10'h8f == idx ? $signed(12'sh477) : $signed(_GEN_142); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_144 = 10'h90 == idx ? $signed(12'sh47f) : $signed(_GEN_143); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_145 = 10'h91 == idx ? $signed(12'sh487) : $signed(_GEN_144); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_146 = 10'h92 == idx ? $signed(12'sh48f) : $signed(_GEN_145); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_147 = 10'h93 == idx ? $signed(12'sh497) : $signed(_GEN_146); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_148 = 10'h94 == idx ? $signed(12'sh49f) : $signed(_GEN_147); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_149 = 10'h95 == idx ? $signed(12'sh4a7) : $signed(_GEN_148); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_150 = 10'h96 == idx ? $signed(12'sh4af) : $signed(_GEN_149); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_151 = 10'h97 == idx ? $signed(12'sh4b7) : $signed(_GEN_150); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_152 = 10'h98 == idx ? $signed(12'sh4bf) : $signed(_GEN_151); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_153 = 10'h99 == idx ? $signed(12'sh4c7) : $signed(_GEN_152); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_154 = 10'h9a == idx ? $signed(12'sh4cf) : $signed(_GEN_153); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_155 = 10'h9b == idx ? $signed(12'sh4d7) : $signed(_GEN_154); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_156 = 10'h9c == idx ? $signed(12'sh4df) : $signed(_GEN_155); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_157 = 10'h9d == idx ? $signed(12'sh4e7) : $signed(_GEN_156); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_158 = 10'h9e == idx ? $signed(12'sh4ef) : $signed(_GEN_157); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_159 = 10'h9f == idx ? $signed(12'sh4f7) : $signed(_GEN_158); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_160 = 10'ha0 == idx ? $signed(12'sh4ff) : $signed(_GEN_159); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_161 = 10'ha1 == idx ? $signed(12'sh507) : $signed(_GEN_160); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_162 = 10'ha2 == idx ? $signed(12'sh50f) : $signed(_GEN_161); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_163 = 10'ha3 == idx ? $signed(12'sh517) : $signed(_GEN_162); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_164 = 10'ha4 == idx ? $signed(12'sh51f) : $signed(_GEN_163); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_165 = 10'ha5 == idx ? $signed(12'sh527) : $signed(_GEN_164); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_166 = 10'ha6 == idx ? $signed(12'sh52f) : $signed(_GEN_165); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_167 = 10'ha7 == idx ? $signed(12'sh537) : $signed(_GEN_166); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_168 = 10'ha8 == idx ? $signed(12'sh53f) : $signed(_GEN_167); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_169 = 10'ha9 == idx ? $signed(12'sh547) : $signed(_GEN_168); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_170 = 10'haa == idx ? $signed(12'sh54f) : $signed(_GEN_169); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_171 = 10'hab == idx ? $signed(12'sh557) : $signed(_GEN_170); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_172 = 10'hac == idx ? $signed(12'sh55f) : $signed(_GEN_171); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_173 = 10'had == idx ? $signed(12'sh567) : $signed(_GEN_172); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_174 = 10'hae == idx ? $signed(12'sh56f) : $signed(_GEN_173); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_175 = 10'haf == idx ? $signed(12'sh577) : $signed(_GEN_174); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_176 = 10'hb0 == idx ? $signed(12'sh57f) : $signed(_GEN_175); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_177 = 10'hb1 == idx ? $signed(12'sh587) : $signed(_GEN_176); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_178 = 10'hb2 == idx ? $signed(12'sh58f) : $signed(_GEN_177); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_179 = 10'hb3 == idx ? $signed(12'sh597) : $signed(_GEN_178); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_180 = 10'hb4 == idx ? $signed(12'sh59f) : $signed(_GEN_179); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_181 = 10'hb5 == idx ? $signed(12'sh5a7) : $signed(_GEN_180); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_182 = 10'hb6 == idx ? $signed(12'sh5af) : $signed(_GEN_181); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_183 = 10'hb7 == idx ? $signed(12'sh5b7) : $signed(_GEN_182); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_184 = 10'hb8 == idx ? $signed(12'sh5bf) : $signed(_GEN_183); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_185 = 10'hb9 == idx ? $signed(12'sh5c7) : $signed(_GEN_184); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_186 = 10'hba == idx ? $signed(12'sh5cf) : $signed(_GEN_185); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_187 = 10'hbb == idx ? $signed(12'sh5d7) : $signed(_GEN_186); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_188 = 10'hbc == idx ? $signed(12'sh5df) : $signed(_GEN_187); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_189 = 10'hbd == idx ? $signed(12'sh5e7) : $signed(_GEN_188); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_190 = 10'hbe == idx ? $signed(12'sh5ef) : $signed(_GEN_189); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_191 = 10'hbf == idx ? $signed(12'sh5f7) : $signed(_GEN_190); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_192 = 10'hc0 == idx ? $signed(12'sh5ff) : $signed(_GEN_191); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_193 = 10'hc1 == idx ? $signed(12'sh607) : $signed(_GEN_192); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_194 = 10'hc2 == idx ? $signed(12'sh60f) : $signed(_GEN_193); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_195 = 10'hc3 == idx ? $signed(12'sh617) : $signed(_GEN_194); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_196 = 10'hc4 == idx ? $signed(12'sh61f) : $signed(_GEN_195); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_197 = 10'hc5 == idx ? $signed(12'sh627) : $signed(_GEN_196); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_198 = 10'hc6 == idx ? $signed(12'sh62f) : $signed(_GEN_197); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_199 = 10'hc7 == idx ? $signed(12'sh637) : $signed(_GEN_198); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_200 = 10'hc8 == idx ? $signed(12'sh63f) : $signed(_GEN_199); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_201 = 10'hc9 == idx ? $signed(12'sh647) : $signed(_GEN_200); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_202 = 10'hca == idx ? $signed(12'sh64f) : $signed(_GEN_201); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_203 = 10'hcb == idx ? $signed(12'sh657) : $signed(_GEN_202); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_204 = 10'hcc == idx ? $signed(12'sh65f) : $signed(_GEN_203); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_205 = 10'hcd == idx ? $signed(12'sh667) : $signed(_GEN_204); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_206 = 10'hce == idx ? $signed(12'sh66f) : $signed(_GEN_205); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_207 = 10'hcf == idx ? $signed(12'sh677) : $signed(_GEN_206); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_208 = 10'hd0 == idx ? $signed(12'sh67f) : $signed(_GEN_207); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_209 = 10'hd1 == idx ? $signed(12'sh687) : $signed(_GEN_208); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_210 = 10'hd2 == idx ? $signed(12'sh68f) : $signed(_GEN_209); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_211 = 10'hd3 == idx ? $signed(12'sh697) : $signed(_GEN_210); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_212 = 10'hd4 == idx ? $signed(12'sh69f) : $signed(_GEN_211); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_213 = 10'hd5 == idx ? $signed(12'sh6a7) : $signed(_GEN_212); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_214 = 10'hd6 == idx ? $signed(12'sh6af) : $signed(_GEN_213); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_215 = 10'hd7 == idx ? $signed(12'sh6b7) : $signed(_GEN_214); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_216 = 10'hd8 == idx ? $signed(12'sh6bf) : $signed(_GEN_215); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_217 = 10'hd9 == idx ? $signed(12'sh6c7) : $signed(_GEN_216); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_218 = 10'hda == idx ? $signed(12'sh6cf) : $signed(_GEN_217); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_219 = 10'hdb == idx ? $signed(12'sh6d7) : $signed(_GEN_218); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_220 = 10'hdc == idx ? $signed(12'sh6df) : $signed(_GEN_219); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_221 = 10'hdd == idx ? $signed(12'sh6e7) : $signed(_GEN_220); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_222 = 10'hde == idx ? $signed(12'sh6ef) : $signed(_GEN_221); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_223 = 10'hdf == idx ? $signed(12'sh6f7) : $signed(_GEN_222); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_224 = 10'he0 == idx ? $signed(12'sh6ff) : $signed(_GEN_223); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_225 = 10'he1 == idx ? $signed(12'sh707) : $signed(_GEN_224); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_226 = 10'he2 == idx ? $signed(12'sh70f) : $signed(_GEN_225); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_227 = 10'he3 == idx ? $signed(12'sh717) : $signed(_GEN_226); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_228 = 10'he4 == idx ? $signed(12'sh71f) : $signed(_GEN_227); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_229 = 10'he5 == idx ? $signed(12'sh727) : $signed(_GEN_228); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_230 = 10'he6 == idx ? $signed(12'sh72f) : $signed(_GEN_229); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_231 = 10'he7 == idx ? $signed(12'sh737) : $signed(_GEN_230); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_232 = 10'he8 == idx ? $signed(12'sh73f) : $signed(_GEN_231); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_233 = 10'he9 == idx ? $signed(12'sh747) : $signed(_GEN_232); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_234 = 10'hea == idx ? $signed(12'sh74f) : $signed(_GEN_233); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_235 = 10'heb == idx ? $signed(12'sh757) : $signed(_GEN_234); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_236 = 10'hec == idx ? $signed(12'sh75f) : $signed(_GEN_235); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_237 = 10'hed == idx ? $signed(12'sh767) : $signed(_GEN_236); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_238 = 10'hee == idx ? $signed(12'sh76f) : $signed(_GEN_237); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_239 = 10'hef == idx ? $signed(12'sh777) : $signed(_GEN_238); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_240 = 10'hf0 == idx ? $signed(12'sh77f) : $signed(_GEN_239); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_241 = 10'hf1 == idx ? $signed(12'sh787) : $signed(_GEN_240); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_242 = 10'hf2 == idx ? $signed(12'sh78f) : $signed(_GEN_241); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_243 = 10'hf3 == idx ? $signed(12'sh797) : $signed(_GEN_242); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_244 = 10'hf4 == idx ? $signed(12'sh79f) : $signed(_GEN_243); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_245 = 10'hf5 == idx ? $signed(12'sh7a7) : $signed(_GEN_244); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_246 = 10'hf6 == idx ? $signed(12'sh7af) : $signed(_GEN_245); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_247 = 10'hf7 == idx ? $signed(12'sh7b7) : $signed(_GEN_246); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_248 = 10'hf8 == idx ? $signed(12'sh7bf) : $signed(_GEN_247); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_249 = 10'hf9 == idx ? $signed(12'sh7c7) : $signed(_GEN_248); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_250 = 10'hfa == idx ? $signed(12'sh7cf) : $signed(_GEN_249); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_251 = 10'hfb == idx ? $signed(12'sh7d7) : $signed(_GEN_250); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_252 = 10'hfc == idx ? $signed(12'sh7df) : $signed(_GEN_251); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_253 = 10'hfd == idx ? $signed(12'sh7e7) : $signed(_GEN_252); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_254 = 10'hfe == idx ? $signed(12'sh7ef) : $signed(_GEN_253); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_255 = 10'hff == idx ? $signed(12'sh7f7) : $signed(_GEN_254); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_256 = 10'h100 == idx ? $signed(12'sh7ff) : $signed(_GEN_255); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_257 = 10'h101 == idx ? $signed(12'sh7f7) : $signed(_GEN_256); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_258 = 10'h102 == idx ? $signed(12'sh7ef) : $signed(_GEN_257); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_259 = 10'h103 == idx ? $signed(12'sh7e7) : $signed(_GEN_258); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_260 = 10'h104 == idx ? $signed(12'sh7df) : $signed(_GEN_259); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_261 = 10'h105 == idx ? $signed(12'sh7d7) : $signed(_GEN_260); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_262 = 10'h106 == idx ? $signed(12'sh7cf) : $signed(_GEN_261); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_263 = 10'h107 == idx ? $signed(12'sh7c7) : $signed(_GEN_262); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_264 = 10'h108 == idx ? $signed(12'sh7bf) : $signed(_GEN_263); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_265 = 10'h109 == idx ? $signed(12'sh7b7) : $signed(_GEN_264); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_266 = 10'h10a == idx ? $signed(12'sh7af) : $signed(_GEN_265); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_267 = 10'h10b == idx ? $signed(12'sh7a7) : $signed(_GEN_266); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_268 = 10'h10c == idx ? $signed(12'sh79f) : $signed(_GEN_267); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_269 = 10'h10d == idx ? $signed(12'sh797) : $signed(_GEN_268); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_270 = 10'h10e == idx ? $signed(12'sh78f) : $signed(_GEN_269); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_271 = 10'h10f == idx ? $signed(12'sh787) : $signed(_GEN_270); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_272 = 10'h110 == idx ? $signed(12'sh77f) : $signed(_GEN_271); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_273 = 10'h111 == idx ? $signed(12'sh777) : $signed(_GEN_272); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_274 = 10'h112 == idx ? $signed(12'sh76f) : $signed(_GEN_273); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_275 = 10'h113 == idx ? $signed(12'sh767) : $signed(_GEN_274); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_276 = 10'h114 == idx ? $signed(12'sh75f) : $signed(_GEN_275); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_277 = 10'h115 == idx ? $signed(12'sh757) : $signed(_GEN_276); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_278 = 10'h116 == idx ? $signed(12'sh74f) : $signed(_GEN_277); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_279 = 10'h117 == idx ? $signed(12'sh747) : $signed(_GEN_278); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_280 = 10'h118 == idx ? $signed(12'sh73f) : $signed(_GEN_279); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_281 = 10'h119 == idx ? $signed(12'sh737) : $signed(_GEN_280); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_282 = 10'h11a == idx ? $signed(12'sh72f) : $signed(_GEN_281); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_283 = 10'h11b == idx ? $signed(12'sh727) : $signed(_GEN_282); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_284 = 10'h11c == idx ? $signed(12'sh71f) : $signed(_GEN_283); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_285 = 10'h11d == idx ? $signed(12'sh717) : $signed(_GEN_284); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_286 = 10'h11e == idx ? $signed(12'sh70f) : $signed(_GEN_285); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_287 = 10'h11f == idx ? $signed(12'sh707) : $signed(_GEN_286); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_288 = 10'h120 == idx ? $signed(12'sh6ff) : $signed(_GEN_287); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_289 = 10'h121 == idx ? $signed(12'sh6f7) : $signed(_GEN_288); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_290 = 10'h122 == idx ? $signed(12'sh6ef) : $signed(_GEN_289); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_291 = 10'h123 == idx ? $signed(12'sh6e7) : $signed(_GEN_290); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_292 = 10'h124 == idx ? $signed(12'sh6df) : $signed(_GEN_291); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_293 = 10'h125 == idx ? $signed(12'sh6d7) : $signed(_GEN_292); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_294 = 10'h126 == idx ? $signed(12'sh6cf) : $signed(_GEN_293); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_295 = 10'h127 == idx ? $signed(12'sh6c7) : $signed(_GEN_294); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_296 = 10'h128 == idx ? $signed(12'sh6bf) : $signed(_GEN_295); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_297 = 10'h129 == idx ? $signed(12'sh6b7) : $signed(_GEN_296); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_298 = 10'h12a == idx ? $signed(12'sh6af) : $signed(_GEN_297); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_299 = 10'h12b == idx ? $signed(12'sh6a7) : $signed(_GEN_298); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_300 = 10'h12c == idx ? $signed(12'sh69f) : $signed(_GEN_299); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_301 = 10'h12d == idx ? $signed(12'sh697) : $signed(_GEN_300); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_302 = 10'h12e == idx ? $signed(12'sh68f) : $signed(_GEN_301); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_303 = 10'h12f == idx ? $signed(12'sh687) : $signed(_GEN_302); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_304 = 10'h130 == idx ? $signed(12'sh67f) : $signed(_GEN_303); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_305 = 10'h131 == idx ? $signed(12'sh677) : $signed(_GEN_304); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_306 = 10'h132 == idx ? $signed(12'sh66f) : $signed(_GEN_305); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_307 = 10'h133 == idx ? $signed(12'sh667) : $signed(_GEN_306); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_308 = 10'h134 == idx ? $signed(12'sh65f) : $signed(_GEN_307); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_309 = 10'h135 == idx ? $signed(12'sh657) : $signed(_GEN_308); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_310 = 10'h136 == idx ? $signed(12'sh64f) : $signed(_GEN_309); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_311 = 10'h137 == idx ? $signed(12'sh647) : $signed(_GEN_310); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_312 = 10'h138 == idx ? $signed(12'sh63f) : $signed(_GEN_311); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_313 = 10'h139 == idx ? $signed(12'sh637) : $signed(_GEN_312); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_314 = 10'h13a == idx ? $signed(12'sh62f) : $signed(_GEN_313); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_315 = 10'h13b == idx ? $signed(12'sh627) : $signed(_GEN_314); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_316 = 10'h13c == idx ? $signed(12'sh61f) : $signed(_GEN_315); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_317 = 10'h13d == idx ? $signed(12'sh617) : $signed(_GEN_316); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_318 = 10'h13e == idx ? $signed(12'sh60f) : $signed(_GEN_317); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_319 = 10'h13f == idx ? $signed(12'sh607) : $signed(_GEN_318); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_320 = 10'h140 == idx ? $signed(12'sh5ff) : $signed(_GEN_319); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_321 = 10'h141 == idx ? $signed(12'sh5f7) : $signed(_GEN_320); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_322 = 10'h142 == idx ? $signed(12'sh5ef) : $signed(_GEN_321); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_323 = 10'h143 == idx ? $signed(12'sh5e7) : $signed(_GEN_322); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_324 = 10'h144 == idx ? $signed(12'sh5df) : $signed(_GEN_323); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_325 = 10'h145 == idx ? $signed(12'sh5d7) : $signed(_GEN_324); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_326 = 10'h146 == idx ? $signed(12'sh5cf) : $signed(_GEN_325); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_327 = 10'h147 == idx ? $signed(12'sh5c7) : $signed(_GEN_326); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_328 = 10'h148 == idx ? $signed(12'sh5bf) : $signed(_GEN_327); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_329 = 10'h149 == idx ? $signed(12'sh5b7) : $signed(_GEN_328); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_330 = 10'h14a == idx ? $signed(12'sh5af) : $signed(_GEN_329); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_331 = 10'h14b == idx ? $signed(12'sh5a7) : $signed(_GEN_330); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_332 = 10'h14c == idx ? $signed(12'sh59f) : $signed(_GEN_331); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_333 = 10'h14d == idx ? $signed(12'sh597) : $signed(_GEN_332); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_334 = 10'h14e == idx ? $signed(12'sh58f) : $signed(_GEN_333); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_335 = 10'h14f == idx ? $signed(12'sh587) : $signed(_GEN_334); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_336 = 10'h150 == idx ? $signed(12'sh57f) : $signed(_GEN_335); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_337 = 10'h151 == idx ? $signed(12'sh577) : $signed(_GEN_336); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_338 = 10'h152 == idx ? $signed(12'sh56f) : $signed(_GEN_337); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_339 = 10'h153 == idx ? $signed(12'sh567) : $signed(_GEN_338); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_340 = 10'h154 == idx ? $signed(12'sh55f) : $signed(_GEN_339); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_341 = 10'h155 == idx ? $signed(12'sh557) : $signed(_GEN_340); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_342 = 10'h156 == idx ? $signed(12'sh54f) : $signed(_GEN_341); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_343 = 10'h157 == idx ? $signed(12'sh547) : $signed(_GEN_342); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_344 = 10'h158 == idx ? $signed(12'sh53f) : $signed(_GEN_343); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_345 = 10'h159 == idx ? $signed(12'sh537) : $signed(_GEN_344); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_346 = 10'h15a == idx ? $signed(12'sh52f) : $signed(_GEN_345); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_347 = 10'h15b == idx ? $signed(12'sh527) : $signed(_GEN_346); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_348 = 10'h15c == idx ? $signed(12'sh51f) : $signed(_GEN_347); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_349 = 10'h15d == idx ? $signed(12'sh517) : $signed(_GEN_348); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_350 = 10'h15e == idx ? $signed(12'sh50f) : $signed(_GEN_349); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_351 = 10'h15f == idx ? $signed(12'sh507) : $signed(_GEN_350); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_352 = 10'h160 == idx ? $signed(12'sh4ff) : $signed(_GEN_351); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_353 = 10'h161 == idx ? $signed(12'sh4f7) : $signed(_GEN_352); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_354 = 10'h162 == idx ? $signed(12'sh4ef) : $signed(_GEN_353); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_355 = 10'h163 == idx ? $signed(12'sh4e7) : $signed(_GEN_354); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_356 = 10'h164 == idx ? $signed(12'sh4df) : $signed(_GEN_355); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_357 = 10'h165 == idx ? $signed(12'sh4d7) : $signed(_GEN_356); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_358 = 10'h166 == idx ? $signed(12'sh4cf) : $signed(_GEN_357); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_359 = 10'h167 == idx ? $signed(12'sh4c7) : $signed(_GEN_358); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_360 = 10'h168 == idx ? $signed(12'sh4bf) : $signed(_GEN_359); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_361 = 10'h169 == idx ? $signed(12'sh4b7) : $signed(_GEN_360); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_362 = 10'h16a == idx ? $signed(12'sh4af) : $signed(_GEN_361); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_363 = 10'h16b == idx ? $signed(12'sh4a7) : $signed(_GEN_362); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_364 = 10'h16c == idx ? $signed(12'sh49f) : $signed(_GEN_363); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_365 = 10'h16d == idx ? $signed(12'sh497) : $signed(_GEN_364); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_366 = 10'h16e == idx ? $signed(12'sh48f) : $signed(_GEN_365); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_367 = 10'h16f == idx ? $signed(12'sh487) : $signed(_GEN_366); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_368 = 10'h170 == idx ? $signed(12'sh47f) : $signed(_GEN_367); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_369 = 10'h171 == idx ? $signed(12'sh477) : $signed(_GEN_368); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_370 = 10'h172 == idx ? $signed(12'sh46f) : $signed(_GEN_369); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_371 = 10'h173 == idx ? $signed(12'sh467) : $signed(_GEN_370); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_372 = 10'h174 == idx ? $signed(12'sh45f) : $signed(_GEN_371); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_373 = 10'h175 == idx ? $signed(12'sh457) : $signed(_GEN_372); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_374 = 10'h176 == idx ? $signed(12'sh44f) : $signed(_GEN_373); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_375 = 10'h177 == idx ? $signed(12'sh447) : $signed(_GEN_374); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_376 = 10'h178 == idx ? $signed(12'sh43f) : $signed(_GEN_375); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_377 = 10'h179 == idx ? $signed(12'sh437) : $signed(_GEN_376); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_378 = 10'h17a == idx ? $signed(12'sh42f) : $signed(_GEN_377); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_379 = 10'h17b == idx ? $signed(12'sh427) : $signed(_GEN_378); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_380 = 10'h17c == idx ? $signed(12'sh41f) : $signed(_GEN_379); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_381 = 10'h17d == idx ? $signed(12'sh417) : $signed(_GEN_380); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_382 = 10'h17e == idx ? $signed(12'sh40f) : $signed(_GEN_381); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_383 = 10'h17f == idx ? $signed(12'sh407) : $signed(_GEN_382); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_384 = 10'h180 == idx ? $signed(12'sh400) : $signed(_GEN_383); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_385 = 10'h181 == idx ? $signed(12'sh3f8) : $signed(_GEN_384); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_386 = 10'h182 == idx ? $signed(12'sh3f0) : $signed(_GEN_385); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_387 = 10'h183 == idx ? $signed(12'sh3e8) : $signed(_GEN_386); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_388 = 10'h184 == idx ? $signed(12'sh3e0) : $signed(_GEN_387); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_389 = 10'h185 == idx ? $signed(12'sh3d8) : $signed(_GEN_388); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_390 = 10'h186 == idx ? $signed(12'sh3d0) : $signed(_GEN_389); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_391 = 10'h187 == idx ? $signed(12'sh3c8) : $signed(_GEN_390); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_392 = 10'h188 == idx ? $signed(12'sh3c0) : $signed(_GEN_391); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_393 = 10'h189 == idx ? $signed(12'sh3b8) : $signed(_GEN_392); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_394 = 10'h18a == idx ? $signed(12'sh3b0) : $signed(_GEN_393); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_395 = 10'h18b == idx ? $signed(12'sh3a8) : $signed(_GEN_394); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_396 = 10'h18c == idx ? $signed(12'sh3a0) : $signed(_GEN_395); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_397 = 10'h18d == idx ? $signed(12'sh398) : $signed(_GEN_396); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_398 = 10'h18e == idx ? $signed(12'sh390) : $signed(_GEN_397); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_399 = 10'h18f == idx ? $signed(12'sh388) : $signed(_GEN_398); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_400 = 10'h190 == idx ? $signed(12'sh380) : $signed(_GEN_399); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_401 = 10'h191 == idx ? $signed(12'sh378) : $signed(_GEN_400); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_402 = 10'h192 == idx ? $signed(12'sh370) : $signed(_GEN_401); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_403 = 10'h193 == idx ? $signed(12'sh368) : $signed(_GEN_402); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_404 = 10'h194 == idx ? $signed(12'sh360) : $signed(_GEN_403); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_405 = 10'h195 == idx ? $signed(12'sh358) : $signed(_GEN_404); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_406 = 10'h196 == idx ? $signed(12'sh350) : $signed(_GEN_405); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_407 = 10'h197 == idx ? $signed(12'sh348) : $signed(_GEN_406); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_408 = 10'h198 == idx ? $signed(12'sh340) : $signed(_GEN_407); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_409 = 10'h199 == idx ? $signed(12'sh338) : $signed(_GEN_408); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_410 = 10'h19a == idx ? $signed(12'sh330) : $signed(_GEN_409); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_411 = 10'h19b == idx ? $signed(12'sh328) : $signed(_GEN_410); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_412 = 10'h19c == idx ? $signed(12'sh320) : $signed(_GEN_411); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_413 = 10'h19d == idx ? $signed(12'sh318) : $signed(_GEN_412); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_414 = 10'h19e == idx ? $signed(12'sh310) : $signed(_GEN_413); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_415 = 10'h19f == idx ? $signed(12'sh308) : $signed(_GEN_414); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_416 = 10'h1a0 == idx ? $signed(12'sh300) : $signed(_GEN_415); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_417 = 10'h1a1 == idx ? $signed(12'sh2f8) : $signed(_GEN_416); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_418 = 10'h1a2 == idx ? $signed(12'sh2f0) : $signed(_GEN_417); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_419 = 10'h1a3 == idx ? $signed(12'sh2e8) : $signed(_GEN_418); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_420 = 10'h1a4 == idx ? $signed(12'sh2e0) : $signed(_GEN_419); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_421 = 10'h1a5 == idx ? $signed(12'sh2d8) : $signed(_GEN_420); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_422 = 10'h1a6 == idx ? $signed(12'sh2d0) : $signed(_GEN_421); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_423 = 10'h1a7 == idx ? $signed(12'sh2c8) : $signed(_GEN_422); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_424 = 10'h1a8 == idx ? $signed(12'sh2c0) : $signed(_GEN_423); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_425 = 10'h1a9 == idx ? $signed(12'sh2b8) : $signed(_GEN_424); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_426 = 10'h1aa == idx ? $signed(12'sh2b0) : $signed(_GEN_425); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_427 = 10'h1ab == idx ? $signed(12'sh2a8) : $signed(_GEN_426); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_428 = 10'h1ac == idx ? $signed(12'sh2a0) : $signed(_GEN_427); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_429 = 10'h1ad == idx ? $signed(12'sh298) : $signed(_GEN_428); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_430 = 10'h1ae == idx ? $signed(12'sh290) : $signed(_GEN_429); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_431 = 10'h1af == idx ? $signed(12'sh288) : $signed(_GEN_430); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_432 = 10'h1b0 == idx ? $signed(12'sh280) : $signed(_GEN_431); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_433 = 10'h1b1 == idx ? $signed(12'sh278) : $signed(_GEN_432); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_434 = 10'h1b2 == idx ? $signed(12'sh270) : $signed(_GEN_433); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_435 = 10'h1b3 == idx ? $signed(12'sh268) : $signed(_GEN_434); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_436 = 10'h1b4 == idx ? $signed(12'sh260) : $signed(_GEN_435); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_437 = 10'h1b5 == idx ? $signed(12'sh258) : $signed(_GEN_436); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_438 = 10'h1b6 == idx ? $signed(12'sh250) : $signed(_GEN_437); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_439 = 10'h1b7 == idx ? $signed(12'sh248) : $signed(_GEN_438); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_440 = 10'h1b8 == idx ? $signed(12'sh240) : $signed(_GEN_439); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_441 = 10'h1b9 == idx ? $signed(12'sh238) : $signed(_GEN_440); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_442 = 10'h1ba == idx ? $signed(12'sh230) : $signed(_GEN_441); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_443 = 10'h1bb == idx ? $signed(12'sh228) : $signed(_GEN_442); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_444 = 10'h1bc == idx ? $signed(12'sh220) : $signed(_GEN_443); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_445 = 10'h1bd == idx ? $signed(12'sh218) : $signed(_GEN_444); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_446 = 10'h1be == idx ? $signed(12'sh210) : $signed(_GEN_445); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_447 = 10'h1bf == idx ? $signed(12'sh208) : $signed(_GEN_446); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_448 = 10'h1c0 == idx ? $signed(12'sh200) : $signed(_GEN_447); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_449 = 10'h1c1 == idx ? $signed(12'sh1f8) : $signed(_GEN_448); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_450 = 10'h1c2 == idx ? $signed(12'sh1f0) : $signed(_GEN_449); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_451 = 10'h1c3 == idx ? $signed(12'sh1e8) : $signed(_GEN_450); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_452 = 10'h1c4 == idx ? $signed(12'sh1e0) : $signed(_GEN_451); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_453 = 10'h1c5 == idx ? $signed(12'sh1d8) : $signed(_GEN_452); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_454 = 10'h1c6 == idx ? $signed(12'sh1d0) : $signed(_GEN_453); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_455 = 10'h1c7 == idx ? $signed(12'sh1c8) : $signed(_GEN_454); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_456 = 10'h1c8 == idx ? $signed(12'sh1c0) : $signed(_GEN_455); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_457 = 10'h1c9 == idx ? $signed(12'sh1b8) : $signed(_GEN_456); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_458 = 10'h1ca == idx ? $signed(12'sh1b0) : $signed(_GEN_457); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_459 = 10'h1cb == idx ? $signed(12'sh1a8) : $signed(_GEN_458); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_460 = 10'h1cc == idx ? $signed(12'sh1a0) : $signed(_GEN_459); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_461 = 10'h1cd == idx ? $signed(12'sh198) : $signed(_GEN_460); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_462 = 10'h1ce == idx ? $signed(12'sh190) : $signed(_GEN_461); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_463 = 10'h1cf == idx ? $signed(12'sh188) : $signed(_GEN_462); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_464 = 10'h1d0 == idx ? $signed(12'sh180) : $signed(_GEN_463); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_465 = 10'h1d1 == idx ? $signed(12'sh178) : $signed(_GEN_464); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_466 = 10'h1d2 == idx ? $signed(12'sh170) : $signed(_GEN_465); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_467 = 10'h1d3 == idx ? $signed(12'sh168) : $signed(_GEN_466); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_468 = 10'h1d4 == idx ? $signed(12'sh160) : $signed(_GEN_467); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_469 = 10'h1d5 == idx ? $signed(12'sh158) : $signed(_GEN_468); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_470 = 10'h1d6 == idx ? $signed(12'sh150) : $signed(_GEN_469); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_471 = 10'h1d7 == idx ? $signed(12'sh148) : $signed(_GEN_470); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_472 = 10'h1d8 == idx ? $signed(12'sh140) : $signed(_GEN_471); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_473 = 10'h1d9 == idx ? $signed(12'sh138) : $signed(_GEN_472); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_474 = 10'h1da == idx ? $signed(12'sh130) : $signed(_GEN_473); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_475 = 10'h1db == idx ? $signed(12'sh128) : $signed(_GEN_474); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_476 = 10'h1dc == idx ? $signed(12'sh120) : $signed(_GEN_475); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_477 = 10'h1dd == idx ? $signed(12'sh118) : $signed(_GEN_476); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_478 = 10'h1de == idx ? $signed(12'sh110) : $signed(_GEN_477); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_479 = 10'h1df == idx ? $signed(12'sh108) : $signed(_GEN_478); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_480 = 10'h1e0 == idx ? $signed(12'sh100) : $signed(_GEN_479); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_481 = 10'h1e1 == idx ? $signed(12'shf8) : $signed(_GEN_480); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_482 = 10'h1e2 == idx ? $signed(12'shf0) : $signed(_GEN_481); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_483 = 10'h1e3 == idx ? $signed(12'she8) : $signed(_GEN_482); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_484 = 10'h1e4 == idx ? $signed(12'she0) : $signed(_GEN_483); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_485 = 10'h1e5 == idx ? $signed(12'shd8) : $signed(_GEN_484); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_486 = 10'h1e6 == idx ? $signed(12'shd0) : $signed(_GEN_485); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_487 = 10'h1e7 == idx ? $signed(12'shc8) : $signed(_GEN_486); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_488 = 10'h1e8 == idx ? $signed(12'shc0) : $signed(_GEN_487); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_489 = 10'h1e9 == idx ? $signed(12'shb8) : $signed(_GEN_488); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_490 = 10'h1ea == idx ? $signed(12'shb0) : $signed(_GEN_489); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_491 = 10'h1eb == idx ? $signed(12'sha8) : $signed(_GEN_490); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_492 = 10'h1ec == idx ? $signed(12'sha0) : $signed(_GEN_491); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_493 = 10'h1ed == idx ? $signed(12'sh98) : $signed(_GEN_492); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_494 = 10'h1ee == idx ? $signed(12'sh90) : $signed(_GEN_493); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_495 = 10'h1ef == idx ? $signed(12'sh88) : $signed(_GEN_494); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_496 = 10'h1f0 == idx ? $signed(12'sh80) : $signed(_GEN_495); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_497 = 10'h1f1 == idx ? $signed(12'sh78) : $signed(_GEN_496); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_498 = 10'h1f2 == idx ? $signed(12'sh70) : $signed(_GEN_497); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_499 = 10'h1f3 == idx ? $signed(12'sh68) : $signed(_GEN_498); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_500 = 10'h1f4 == idx ? $signed(12'sh60) : $signed(_GEN_499); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_501 = 10'h1f5 == idx ? $signed(12'sh58) : $signed(_GEN_500); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_502 = 10'h1f6 == idx ? $signed(12'sh50) : $signed(_GEN_501); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_503 = 10'h1f7 == idx ? $signed(12'sh48) : $signed(_GEN_502); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_504 = 10'h1f8 == idx ? $signed(12'sh40) : $signed(_GEN_503); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_505 = 10'h1f9 == idx ? $signed(12'sh38) : $signed(_GEN_504); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_506 = 10'h1fa == idx ? $signed(12'sh30) : $signed(_GEN_505); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_507 = 10'h1fb == idx ? $signed(12'sh28) : $signed(_GEN_506); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_508 = 10'h1fc == idx ? $signed(12'sh20) : $signed(_GEN_507); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_509 = 10'h1fd == idx ? $signed(12'sh18) : $signed(_GEN_508); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_510 = 10'h1fe == idx ? $signed(12'sh10) : $signed(_GEN_509); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_511 = 10'h1ff == idx ? $signed(12'sh8) : $signed(_GEN_510); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_512 = 10'h200 == idx ? $signed(12'sh0) : $signed(_GEN_511); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_513 = 10'h201 == idx ? $signed(-12'sh8) : $signed(_GEN_512); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_514 = 10'h202 == idx ? $signed(-12'sh10) : $signed(_GEN_513); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_515 = 10'h203 == idx ? $signed(-12'sh18) : $signed(_GEN_514); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_516 = 10'h204 == idx ? $signed(-12'sh20) : $signed(_GEN_515); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_517 = 10'h205 == idx ? $signed(-12'sh28) : $signed(_GEN_516); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_518 = 10'h206 == idx ? $signed(-12'sh30) : $signed(_GEN_517); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_519 = 10'h207 == idx ? $signed(-12'sh38) : $signed(_GEN_518); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_520 = 10'h208 == idx ? $signed(-12'sh40) : $signed(_GEN_519); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_521 = 10'h209 == idx ? $signed(-12'sh48) : $signed(_GEN_520); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_522 = 10'h20a == idx ? $signed(-12'sh50) : $signed(_GEN_521); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_523 = 10'h20b == idx ? $signed(-12'sh58) : $signed(_GEN_522); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_524 = 10'h20c == idx ? $signed(-12'sh60) : $signed(_GEN_523); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_525 = 10'h20d == idx ? $signed(-12'sh68) : $signed(_GEN_524); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_526 = 10'h20e == idx ? $signed(-12'sh70) : $signed(_GEN_525); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_527 = 10'h20f == idx ? $signed(-12'sh78) : $signed(_GEN_526); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_528 = 10'h210 == idx ? $signed(-12'sh80) : $signed(_GEN_527); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_529 = 10'h211 == idx ? $signed(-12'sh88) : $signed(_GEN_528); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_530 = 10'h212 == idx ? $signed(-12'sh90) : $signed(_GEN_529); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_531 = 10'h213 == idx ? $signed(-12'sh98) : $signed(_GEN_530); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_532 = 10'h214 == idx ? $signed(-12'sha0) : $signed(_GEN_531); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_533 = 10'h215 == idx ? $signed(-12'sha8) : $signed(_GEN_532); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_534 = 10'h216 == idx ? $signed(-12'shb0) : $signed(_GEN_533); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_535 = 10'h217 == idx ? $signed(-12'shb8) : $signed(_GEN_534); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_536 = 10'h218 == idx ? $signed(-12'shc0) : $signed(_GEN_535); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_537 = 10'h219 == idx ? $signed(-12'shc8) : $signed(_GEN_536); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_538 = 10'h21a == idx ? $signed(-12'shd0) : $signed(_GEN_537); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_539 = 10'h21b == idx ? $signed(-12'shd8) : $signed(_GEN_538); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_540 = 10'h21c == idx ? $signed(-12'she0) : $signed(_GEN_539); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_541 = 10'h21d == idx ? $signed(-12'she8) : $signed(_GEN_540); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_542 = 10'h21e == idx ? $signed(-12'shf0) : $signed(_GEN_541); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_543 = 10'h21f == idx ? $signed(-12'shf8) : $signed(_GEN_542); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_544 = 10'h220 == idx ? $signed(-12'sh100) : $signed(_GEN_543); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_545 = 10'h221 == idx ? $signed(-12'sh108) : $signed(_GEN_544); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_546 = 10'h222 == idx ? $signed(-12'sh110) : $signed(_GEN_545); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_547 = 10'h223 == idx ? $signed(-12'sh118) : $signed(_GEN_546); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_548 = 10'h224 == idx ? $signed(-12'sh120) : $signed(_GEN_547); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_549 = 10'h225 == idx ? $signed(-12'sh128) : $signed(_GEN_548); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_550 = 10'h226 == idx ? $signed(-12'sh130) : $signed(_GEN_549); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_551 = 10'h227 == idx ? $signed(-12'sh138) : $signed(_GEN_550); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_552 = 10'h228 == idx ? $signed(-12'sh140) : $signed(_GEN_551); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_553 = 10'h229 == idx ? $signed(-12'sh148) : $signed(_GEN_552); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_554 = 10'h22a == idx ? $signed(-12'sh150) : $signed(_GEN_553); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_555 = 10'h22b == idx ? $signed(-12'sh158) : $signed(_GEN_554); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_556 = 10'h22c == idx ? $signed(-12'sh160) : $signed(_GEN_555); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_557 = 10'h22d == idx ? $signed(-12'sh168) : $signed(_GEN_556); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_558 = 10'h22e == idx ? $signed(-12'sh170) : $signed(_GEN_557); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_559 = 10'h22f == idx ? $signed(-12'sh178) : $signed(_GEN_558); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_560 = 10'h230 == idx ? $signed(-12'sh180) : $signed(_GEN_559); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_561 = 10'h231 == idx ? $signed(-12'sh188) : $signed(_GEN_560); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_562 = 10'h232 == idx ? $signed(-12'sh190) : $signed(_GEN_561); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_563 = 10'h233 == idx ? $signed(-12'sh198) : $signed(_GEN_562); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_564 = 10'h234 == idx ? $signed(-12'sh1a0) : $signed(_GEN_563); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_565 = 10'h235 == idx ? $signed(-12'sh1a8) : $signed(_GEN_564); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_566 = 10'h236 == idx ? $signed(-12'sh1b0) : $signed(_GEN_565); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_567 = 10'h237 == idx ? $signed(-12'sh1b8) : $signed(_GEN_566); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_568 = 10'h238 == idx ? $signed(-12'sh1c0) : $signed(_GEN_567); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_569 = 10'h239 == idx ? $signed(-12'sh1c8) : $signed(_GEN_568); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_570 = 10'h23a == idx ? $signed(-12'sh1d0) : $signed(_GEN_569); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_571 = 10'h23b == idx ? $signed(-12'sh1d8) : $signed(_GEN_570); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_572 = 10'h23c == idx ? $signed(-12'sh1e0) : $signed(_GEN_571); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_573 = 10'h23d == idx ? $signed(-12'sh1e8) : $signed(_GEN_572); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_574 = 10'h23e == idx ? $signed(-12'sh1f0) : $signed(_GEN_573); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_575 = 10'h23f == idx ? $signed(-12'sh1f8) : $signed(_GEN_574); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_576 = 10'h240 == idx ? $signed(-12'sh200) : $signed(_GEN_575); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_577 = 10'h241 == idx ? $signed(-12'sh208) : $signed(_GEN_576); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_578 = 10'h242 == idx ? $signed(-12'sh210) : $signed(_GEN_577); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_579 = 10'h243 == idx ? $signed(-12'sh218) : $signed(_GEN_578); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_580 = 10'h244 == idx ? $signed(-12'sh220) : $signed(_GEN_579); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_581 = 10'h245 == idx ? $signed(-12'sh228) : $signed(_GEN_580); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_582 = 10'h246 == idx ? $signed(-12'sh230) : $signed(_GEN_581); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_583 = 10'h247 == idx ? $signed(-12'sh238) : $signed(_GEN_582); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_584 = 10'h248 == idx ? $signed(-12'sh240) : $signed(_GEN_583); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_585 = 10'h249 == idx ? $signed(-12'sh248) : $signed(_GEN_584); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_586 = 10'h24a == idx ? $signed(-12'sh250) : $signed(_GEN_585); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_587 = 10'h24b == idx ? $signed(-12'sh258) : $signed(_GEN_586); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_588 = 10'h24c == idx ? $signed(-12'sh260) : $signed(_GEN_587); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_589 = 10'h24d == idx ? $signed(-12'sh268) : $signed(_GEN_588); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_590 = 10'h24e == idx ? $signed(-12'sh270) : $signed(_GEN_589); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_591 = 10'h24f == idx ? $signed(-12'sh278) : $signed(_GEN_590); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_592 = 10'h250 == idx ? $signed(-12'sh280) : $signed(_GEN_591); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_593 = 10'h251 == idx ? $signed(-12'sh288) : $signed(_GEN_592); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_594 = 10'h252 == idx ? $signed(-12'sh290) : $signed(_GEN_593); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_595 = 10'h253 == idx ? $signed(-12'sh298) : $signed(_GEN_594); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_596 = 10'h254 == idx ? $signed(-12'sh2a0) : $signed(_GEN_595); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_597 = 10'h255 == idx ? $signed(-12'sh2a8) : $signed(_GEN_596); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_598 = 10'h256 == idx ? $signed(-12'sh2b0) : $signed(_GEN_597); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_599 = 10'h257 == idx ? $signed(-12'sh2b8) : $signed(_GEN_598); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_600 = 10'h258 == idx ? $signed(-12'sh2c0) : $signed(_GEN_599); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_601 = 10'h259 == idx ? $signed(-12'sh2c8) : $signed(_GEN_600); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_602 = 10'h25a == idx ? $signed(-12'sh2d0) : $signed(_GEN_601); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_603 = 10'h25b == idx ? $signed(-12'sh2d8) : $signed(_GEN_602); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_604 = 10'h25c == idx ? $signed(-12'sh2e0) : $signed(_GEN_603); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_605 = 10'h25d == idx ? $signed(-12'sh2e8) : $signed(_GEN_604); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_606 = 10'h25e == idx ? $signed(-12'sh2f0) : $signed(_GEN_605); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_607 = 10'h25f == idx ? $signed(-12'sh2f8) : $signed(_GEN_606); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_608 = 10'h260 == idx ? $signed(-12'sh300) : $signed(_GEN_607); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_609 = 10'h261 == idx ? $signed(-12'sh308) : $signed(_GEN_608); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_610 = 10'h262 == idx ? $signed(-12'sh310) : $signed(_GEN_609); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_611 = 10'h263 == idx ? $signed(-12'sh318) : $signed(_GEN_610); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_612 = 10'h264 == idx ? $signed(-12'sh320) : $signed(_GEN_611); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_613 = 10'h265 == idx ? $signed(-12'sh328) : $signed(_GEN_612); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_614 = 10'h266 == idx ? $signed(-12'sh330) : $signed(_GEN_613); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_615 = 10'h267 == idx ? $signed(-12'sh338) : $signed(_GEN_614); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_616 = 10'h268 == idx ? $signed(-12'sh340) : $signed(_GEN_615); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_617 = 10'h269 == idx ? $signed(-12'sh348) : $signed(_GEN_616); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_618 = 10'h26a == idx ? $signed(-12'sh350) : $signed(_GEN_617); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_619 = 10'h26b == idx ? $signed(-12'sh358) : $signed(_GEN_618); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_620 = 10'h26c == idx ? $signed(-12'sh360) : $signed(_GEN_619); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_621 = 10'h26d == idx ? $signed(-12'sh368) : $signed(_GEN_620); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_622 = 10'h26e == idx ? $signed(-12'sh370) : $signed(_GEN_621); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_623 = 10'h26f == idx ? $signed(-12'sh378) : $signed(_GEN_622); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_624 = 10'h270 == idx ? $signed(-12'sh380) : $signed(_GEN_623); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_625 = 10'h271 == idx ? $signed(-12'sh388) : $signed(_GEN_624); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_626 = 10'h272 == idx ? $signed(-12'sh390) : $signed(_GEN_625); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_627 = 10'h273 == idx ? $signed(-12'sh398) : $signed(_GEN_626); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_628 = 10'h274 == idx ? $signed(-12'sh3a0) : $signed(_GEN_627); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_629 = 10'h275 == idx ? $signed(-12'sh3a8) : $signed(_GEN_628); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_630 = 10'h276 == idx ? $signed(-12'sh3b0) : $signed(_GEN_629); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_631 = 10'h277 == idx ? $signed(-12'sh3b8) : $signed(_GEN_630); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_632 = 10'h278 == idx ? $signed(-12'sh3c0) : $signed(_GEN_631); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_633 = 10'h279 == idx ? $signed(-12'sh3c8) : $signed(_GEN_632); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_634 = 10'h27a == idx ? $signed(-12'sh3d0) : $signed(_GEN_633); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_635 = 10'h27b == idx ? $signed(-12'sh3d8) : $signed(_GEN_634); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_636 = 10'h27c == idx ? $signed(-12'sh3e0) : $signed(_GEN_635); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_637 = 10'h27d == idx ? $signed(-12'sh3e8) : $signed(_GEN_636); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_638 = 10'h27e == idx ? $signed(-12'sh3f0) : $signed(_GEN_637); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_639 = 10'h27f == idx ? $signed(-12'sh3f8) : $signed(_GEN_638); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_640 = 10'h280 == idx ? $signed(-12'sh3ff) : $signed(_GEN_639); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_641 = 10'h281 == idx ? $signed(-12'sh407) : $signed(_GEN_640); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_642 = 10'h282 == idx ? $signed(-12'sh40f) : $signed(_GEN_641); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_643 = 10'h283 == idx ? $signed(-12'sh417) : $signed(_GEN_642); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_644 = 10'h284 == idx ? $signed(-12'sh41f) : $signed(_GEN_643); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_645 = 10'h285 == idx ? $signed(-12'sh427) : $signed(_GEN_644); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_646 = 10'h286 == idx ? $signed(-12'sh42f) : $signed(_GEN_645); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_647 = 10'h287 == idx ? $signed(-12'sh437) : $signed(_GEN_646); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_648 = 10'h288 == idx ? $signed(-12'sh43f) : $signed(_GEN_647); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_649 = 10'h289 == idx ? $signed(-12'sh447) : $signed(_GEN_648); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_650 = 10'h28a == idx ? $signed(-12'sh44f) : $signed(_GEN_649); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_651 = 10'h28b == idx ? $signed(-12'sh457) : $signed(_GEN_650); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_652 = 10'h28c == idx ? $signed(-12'sh45f) : $signed(_GEN_651); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_653 = 10'h28d == idx ? $signed(-12'sh467) : $signed(_GEN_652); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_654 = 10'h28e == idx ? $signed(-12'sh46f) : $signed(_GEN_653); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_655 = 10'h28f == idx ? $signed(-12'sh477) : $signed(_GEN_654); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_656 = 10'h290 == idx ? $signed(-12'sh47f) : $signed(_GEN_655); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_657 = 10'h291 == idx ? $signed(-12'sh487) : $signed(_GEN_656); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_658 = 10'h292 == idx ? $signed(-12'sh48f) : $signed(_GEN_657); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_659 = 10'h293 == idx ? $signed(-12'sh497) : $signed(_GEN_658); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_660 = 10'h294 == idx ? $signed(-12'sh49f) : $signed(_GEN_659); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_661 = 10'h295 == idx ? $signed(-12'sh4a7) : $signed(_GEN_660); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_662 = 10'h296 == idx ? $signed(-12'sh4af) : $signed(_GEN_661); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_663 = 10'h297 == idx ? $signed(-12'sh4b7) : $signed(_GEN_662); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_664 = 10'h298 == idx ? $signed(-12'sh4bf) : $signed(_GEN_663); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_665 = 10'h299 == idx ? $signed(-12'sh4c7) : $signed(_GEN_664); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_666 = 10'h29a == idx ? $signed(-12'sh4cf) : $signed(_GEN_665); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_667 = 10'h29b == idx ? $signed(-12'sh4d7) : $signed(_GEN_666); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_668 = 10'h29c == idx ? $signed(-12'sh4df) : $signed(_GEN_667); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_669 = 10'h29d == idx ? $signed(-12'sh4e7) : $signed(_GEN_668); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_670 = 10'h29e == idx ? $signed(-12'sh4ef) : $signed(_GEN_669); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_671 = 10'h29f == idx ? $signed(-12'sh4f7) : $signed(_GEN_670); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_672 = 10'h2a0 == idx ? $signed(-12'sh4ff) : $signed(_GEN_671); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_673 = 10'h2a1 == idx ? $signed(-12'sh507) : $signed(_GEN_672); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_674 = 10'h2a2 == idx ? $signed(-12'sh50f) : $signed(_GEN_673); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_675 = 10'h2a3 == idx ? $signed(-12'sh517) : $signed(_GEN_674); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_676 = 10'h2a4 == idx ? $signed(-12'sh51f) : $signed(_GEN_675); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_677 = 10'h2a5 == idx ? $signed(-12'sh527) : $signed(_GEN_676); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_678 = 10'h2a6 == idx ? $signed(-12'sh52f) : $signed(_GEN_677); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_679 = 10'h2a7 == idx ? $signed(-12'sh537) : $signed(_GEN_678); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_680 = 10'h2a8 == idx ? $signed(-12'sh53f) : $signed(_GEN_679); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_681 = 10'h2a9 == idx ? $signed(-12'sh547) : $signed(_GEN_680); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_682 = 10'h2aa == idx ? $signed(-12'sh54f) : $signed(_GEN_681); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_683 = 10'h2ab == idx ? $signed(-12'sh557) : $signed(_GEN_682); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_684 = 10'h2ac == idx ? $signed(-12'sh55f) : $signed(_GEN_683); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_685 = 10'h2ad == idx ? $signed(-12'sh567) : $signed(_GEN_684); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_686 = 10'h2ae == idx ? $signed(-12'sh56f) : $signed(_GEN_685); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_687 = 10'h2af == idx ? $signed(-12'sh577) : $signed(_GEN_686); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_688 = 10'h2b0 == idx ? $signed(-12'sh57f) : $signed(_GEN_687); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_689 = 10'h2b1 == idx ? $signed(-12'sh587) : $signed(_GEN_688); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_690 = 10'h2b2 == idx ? $signed(-12'sh58f) : $signed(_GEN_689); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_691 = 10'h2b3 == idx ? $signed(-12'sh597) : $signed(_GEN_690); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_692 = 10'h2b4 == idx ? $signed(-12'sh59f) : $signed(_GEN_691); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_693 = 10'h2b5 == idx ? $signed(-12'sh5a7) : $signed(_GEN_692); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_694 = 10'h2b6 == idx ? $signed(-12'sh5af) : $signed(_GEN_693); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_695 = 10'h2b7 == idx ? $signed(-12'sh5b7) : $signed(_GEN_694); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_696 = 10'h2b8 == idx ? $signed(-12'sh5bf) : $signed(_GEN_695); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_697 = 10'h2b9 == idx ? $signed(-12'sh5c7) : $signed(_GEN_696); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_698 = 10'h2ba == idx ? $signed(-12'sh5cf) : $signed(_GEN_697); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_699 = 10'h2bb == idx ? $signed(-12'sh5d7) : $signed(_GEN_698); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_700 = 10'h2bc == idx ? $signed(-12'sh5df) : $signed(_GEN_699); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_701 = 10'h2bd == idx ? $signed(-12'sh5e7) : $signed(_GEN_700); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_702 = 10'h2be == idx ? $signed(-12'sh5ef) : $signed(_GEN_701); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_703 = 10'h2bf == idx ? $signed(-12'sh5f7) : $signed(_GEN_702); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_704 = 10'h2c0 == idx ? $signed(-12'sh5ff) : $signed(_GEN_703); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_705 = 10'h2c1 == idx ? $signed(-12'sh607) : $signed(_GEN_704); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_706 = 10'h2c2 == idx ? $signed(-12'sh60f) : $signed(_GEN_705); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_707 = 10'h2c3 == idx ? $signed(-12'sh617) : $signed(_GEN_706); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_708 = 10'h2c4 == idx ? $signed(-12'sh61f) : $signed(_GEN_707); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_709 = 10'h2c5 == idx ? $signed(-12'sh627) : $signed(_GEN_708); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_710 = 10'h2c6 == idx ? $signed(-12'sh62f) : $signed(_GEN_709); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_711 = 10'h2c7 == idx ? $signed(-12'sh637) : $signed(_GEN_710); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_712 = 10'h2c8 == idx ? $signed(-12'sh63f) : $signed(_GEN_711); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_713 = 10'h2c9 == idx ? $signed(-12'sh647) : $signed(_GEN_712); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_714 = 10'h2ca == idx ? $signed(-12'sh64f) : $signed(_GEN_713); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_715 = 10'h2cb == idx ? $signed(-12'sh657) : $signed(_GEN_714); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_716 = 10'h2cc == idx ? $signed(-12'sh65f) : $signed(_GEN_715); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_717 = 10'h2cd == idx ? $signed(-12'sh667) : $signed(_GEN_716); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_718 = 10'h2ce == idx ? $signed(-12'sh66f) : $signed(_GEN_717); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_719 = 10'h2cf == idx ? $signed(-12'sh677) : $signed(_GEN_718); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_720 = 10'h2d0 == idx ? $signed(-12'sh67f) : $signed(_GEN_719); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_721 = 10'h2d1 == idx ? $signed(-12'sh687) : $signed(_GEN_720); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_722 = 10'h2d2 == idx ? $signed(-12'sh68f) : $signed(_GEN_721); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_723 = 10'h2d3 == idx ? $signed(-12'sh697) : $signed(_GEN_722); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_724 = 10'h2d4 == idx ? $signed(-12'sh69f) : $signed(_GEN_723); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_725 = 10'h2d5 == idx ? $signed(-12'sh6a7) : $signed(_GEN_724); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_726 = 10'h2d6 == idx ? $signed(-12'sh6af) : $signed(_GEN_725); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_727 = 10'h2d7 == idx ? $signed(-12'sh6b7) : $signed(_GEN_726); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_728 = 10'h2d8 == idx ? $signed(-12'sh6bf) : $signed(_GEN_727); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_729 = 10'h2d9 == idx ? $signed(-12'sh6c7) : $signed(_GEN_728); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_730 = 10'h2da == idx ? $signed(-12'sh6cf) : $signed(_GEN_729); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_731 = 10'h2db == idx ? $signed(-12'sh6d7) : $signed(_GEN_730); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_732 = 10'h2dc == idx ? $signed(-12'sh6df) : $signed(_GEN_731); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_733 = 10'h2dd == idx ? $signed(-12'sh6e7) : $signed(_GEN_732); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_734 = 10'h2de == idx ? $signed(-12'sh6ef) : $signed(_GEN_733); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_735 = 10'h2df == idx ? $signed(-12'sh6f7) : $signed(_GEN_734); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_736 = 10'h2e0 == idx ? $signed(-12'sh6ff) : $signed(_GEN_735); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_737 = 10'h2e1 == idx ? $signed(-12'sh707) : $signed(_GEN_736); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_738 = 10'h2e2 == idx ? $signed(-12'sh70f) : $signed(_GEN_737); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_739 = 10'h2e3 == idx ? $signed(-12'sh717) : $signed(_GEN_738); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_740 = 10'h2e4 == idx ? $signed(-12'sh71f) : $signed(_GEN_739); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_741 = 10'h2e5 == idx ? $signed(-12'sh727) : $signed(_GEN_740); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_742 = 10'h2e6 == idx ? $signed(-12'sh72f) : $signed(_GEN_741); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_743 = 10'h2e7 == idx ? $signed(-12'sh737) : $signed(_GEN_742); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_744 = 10'h2e8 == idx ? $signed(-12'sh73f) : $signed(_GEN_743); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_745 = 10'h2e9 == idx ? $signed(-12'sh747) : $signed(_GEN_744); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_746 = 10'h2ea == idx ? $signed(-12'sh74f) : $signed(_GEN_745); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_747 = 10'h2eb == idx ? $signed(-12'sh757) : $signed(_GEN_746); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_748 = 10'h2ec == idx ? $signed(-12'sh75f) : $signed(_GEN_747); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_749 = 10'h2ed == idx ? $signed(-12'sh767) : $signed(_GEN_748); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_750 = 10'h2ee == idx ? $signed(-12'sh76f) : $signed(_GEN_749); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_751 = 10'h2ef == idx ? $signed(-12'sh777) : $signed(_GEN_750); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_752 = 10'h2f0 == idx ? $signed(-12'sh77f) : $signed(_GEN_751); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_753 = 10'h2f1 == idx ? $signed(-12'sh787) : $signed(_GEN_752); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_754 = 10'h2f2 == idx ? $signed(-12'sh78f) : $signed(_GEN_753); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_755 = 10'h2f3 == idx ? $signed(-12'sh797) : $signed(_GEN_754); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_756 = 10'h2f4 == idx ? $signed(-12'sh79f) : $signed(_GEN_755); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_757 = 10'h2f5 == idx ? $signed(-12'sh7a7) : $signed(_GEN_756); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_758 = 10'h2f6 == idx ? $signed(-12'sh7af) : $signed(_GEN_757); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_759 = 10'h2f7 == idx ? $signed(-12'sh7b7) : $signed(_GEN_758); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_760 = 10'h2f8 == idx ? $signed(-12'sh7bf) : $signed(_GEN_759); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_761 = 10'h2f9 == idx ? $signed(-12'sh7c7) : $signed(_GEN_760); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_762 = 10'h2fa == idx ? $signed(-12'sh7cf) : $signed(_GEN_761); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_763 = 10'h2fb == idx ? $signed(-12'sh7d7) : $signed(_GEN_762); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_764 = 10'h2fc == idx ? $signed(-12'sh7df) : $signed(_GEN_763); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_765 = 10'h2fd == idx ? $signed(-12'sh7e7) : $signed(_GEN_764); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_766 = 10'h2fe == idx ? $signed(-12'sh7ef) : $signed(_GEN_765); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_767 = 10'h2ff == idx ? $signed(-12'sh7f7) : $signed(_GEN_766); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_768 = 10'h300 == idx ? $signed(-12'sh7ff) : $signed(_GEN_767); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_769 = 10'h301 == idx ? $signed(-12'sh7f7) : $signed(_GEN_768); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_770 = 10'h302 == idx ? $signed(-12'sh7ef) : $signed(_GEN_769); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_771 = 10'h303 == idx ? $signed(-12'sh7e7) : $signed(_GEN_770); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_772 = 10'h304 == idx ? $signed(-12'sh7df) : $signed(_GEN_771); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_773 = 10'h305 == idx ? $signed(-12'sh7d7) : $signed(_GEN_772); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_774 = 10'h306 == idx ? $signed(-12'sh7cf) : $signed(_GEN_773); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_775 = 10'h307 == idx ? $signed(-12'sh7c7) : $signed(_GEN_774); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_776 = 10'h308 == idx ? $signed(-12'sh7bf) : $signed(_GEN_775); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_777 = 10'h309 == idx ? $signed(-12'sh7b7) : $signed(_GEN_776); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_778 = 10'h30a == idx ? $signed(-12'sh7af) : $signed(_GEN_777); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_779 = 10'h30b == idx ? $signed(-12'sh7a7) : $signed(_GEN_778); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_780 = 10'h30c == idx ? $signed(-12'sh79f) : $signed(_GEN_779); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_781 = 10'h30d == idx ? $signed(-12'sh797) : $signed(_GEN_780); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_782 = 10'h30e == idx ? $signed(-12'sh78f) : $signed(_GEN_781); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_783 = 10'h30f == idx ? $signed(-12'sh787) : $signed(_GEN_782); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_784 = 10'h310 == idx ? $signed(-12'sh77f) : $signed(_GEN_783); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_785 = 10'h311 == idx ? $signed(-12'sh777) : $signed(_GEN_784); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_786 = 10'h312 == idx ? $signed(-12'sh76f) : $signed(_GEN_785); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_787 = 10'h313 == idx ? $signed(-12'sh767) : $signed(_GEN_786); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_788 = 10'h314 == idx ? $signed(-12'sh75f) : $signed(_GEN_787); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_789 = 10'h315 == idx ? $signed(-12'sh757) : $signed(_GEN_788); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_790 = 10'h316 == idx ? $signed(-12'sh74f) : $signed(_GEN_789); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_791 = 10'h317 == idx ? $signed(-12'sh747) : $signed(_GEN_790); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_792 = 10'h318 == idx ? $signed(-12'sh73f) : $signed(_GEN_791); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_793 = 10'h319 == idx ? $signed(-12'sh737) : $signed(_GEN_792); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_794 = 10'h31a == idx ? $signed(-12'sh72f) : $signed(_GEN_793); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_795 = 10'h31b == idx ? $signed(-12'sh727) : $signed(_GEN_794); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_796 = 10'h31c == idx ? $signed(-12'sh71f) : $signed(_GEN_795); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_797 = 10'h31d == idx ? $signed(-12'sh717) : $signed(_GEN_796); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_798 = 10'h31e == idx ? $signed(-12'sh70f) : $signed(_GEN_797); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_799 = 10'h31f == idx ? $signed(-12'sh707) : $signed(_GEN_798); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_800 = 10'h320 == idx ? $signed(-12'sh6ff) : $signed(_GEN_799); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_801 = 10'h321 == idx ? $signed(-12'sh6f7) : $signed(_GEN_800); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_802 = 10'h322 == idx ? $signed(-12'sh6ef) : $signed(_GEN_801); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_803 = 10'h323 == idx ? $signed(-12'sh6e7) : $signed(_GEN_802); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_804 = 10'h324 == idx ? $signed(-12'sh6df) : $signed(_GEN_803); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_805 = 10'h325 == idx ? $signed(-12'sh6d7) : $signed(_GEN_804); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_806 = 10'h326 == idx ? $signed(-12'sh6cf) : $signed(_GEN_805); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_807 = 10'h327 == idx ? $signed(-12'sh6c7) : $signed(_GEN_806); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_808 = 10'h328 == idx ? $signed(-12'sh6bf) : $signed(_GEN_807); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_809 = 10'h329 == idx ? $signed(-12'sh6b7) : $signed(_GEN_808); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_810 = 10'h32a == idx ? $signed(-12'sh6af) : $signed(_GEN_809); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_811 = 10'h32b == idx ? $signed(-12'sh6a7) : $signed(_GEN_810); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_812 = 10'h32c == idx ? $signed(-12'sh69f) : $signed(_GEN_811); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_813 = 10'h32d == idx ? $signed(-12'sh697) : $signed(_GEN_812); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_814 = 10'h32e == idx ? $signed(-12'sh68f) : $signed(_GEN_813); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_815 = 10'h32f == idx ? $signed(-12'sh687) : $signed(_GEN_814); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_816 = 10'h330 == idx ? $signed(-12'sh67f) : $signed(_GEN_815); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_817 = 10'h331 == idx ? $signed(-12'sh677) : $signed(_GEN_816); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_818 = 10'h332 == idx ? $signed(-12'sh66f) : $signed(_GEN_817); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_819 = 10'h333 == idx ? $signed(-12'sh667) : $signed(_GEN_818); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_820 = 10'h334 == idx ? $signed(-12'sh65f) : $signed(_GEN_819); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_821 = 10'h335 == idx ? $signed(-12'sh657) : $signed(_GEN_820); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_822 = 10'h336 == idx ? $signed(-12'sh64f) : $signed(_GEN_821); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_823 = 10'h337 == idx ? $signed(-12'sh647) : $signed(_GEN_822); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_824 = 10'h338 == idx ? $signed(-12'sh63f) : $signed(_GEN_823); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_825 = 10'h339 == idx ? $signed(-12'sh637) : $signed(_GEN_824); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_826 = 10'h33a == idx ? $signed(-12'sh62f) : $signed(_GEN_825); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_827 = 10'h33b == idx ? $signed(-12'sh627) : $signed(_GEN_826); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_828 = 10'h33c == idx ? $signed(-12'sh61f) : $signed(_GEN_827); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_829 = 10'h33d == idx ? $signed(-12'sh617) : $signed(_GEN_828); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_830 = 10'h33e == idx ? $signed(-12'sh60f) : $signed(_GEN_829); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_831 = 10'h33f == idx ? $signed(-12'sh607) : $signed(_GEN_830); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_832 = 10'h340 == idx ? $signed(-12'sh5ff) : $signed(_GEN_831); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_833 = 10'h341 == idx ? $signed(-12'sh5f7) : $signed(_GEN_832); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_834 = 10'h342 == idx ? $signed(-12'sh5ef) : $signed(_GEN_833); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_835 = 10'h343 == idx ? $signed(-12'sh5e7) : $signed(_GEN_834); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_836 = 10'h344 == idx ? $signed(-12'sh5df) : $signed(_GEN_835); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_837 = 10'h345 == idx ? $signed(-12'sh5d7) : $signed(_GEN_836); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_838 = 10'h346 == idx ? $signed(-12'sh5cf) : $signed(_GEN_837); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_839 = 10'h347 == idx ? $signed(-12'sh5c7) : $signed(_GEN_838); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_840 = 10'h348 == idx ? $signed(-12'sh5bf) : $signed(_GEN_839); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_841 = 10'h349 == idx ? $signed(-12'sh5b7) : $signed(_GEN_840); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_842 = 10'h34a == idx ? $signed(-12'sh5af) : $signed(_GEN_841); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_843 = 10'h34b == idx ? $signed(-12'sh5a7) : $signed(_GEN_842); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_844 = 10'h34c == idx ? $signed(-12'sh59f) : $signed(_GEN_843); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_845 = 10'h34d == idx ? $signed(-12'sh597) : $signed(_GEN_844); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_846 = 10'h34e == idx ? $signed(-12'sh58f) : $signed(_GEN_845); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_847 = 10'h34f == idx ? $signed(-12'sh587) : $signed(_GEN_846); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_848 = 10'h350 == idx ? $signed(-12'sh57f) : $signed(_GEN_847); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_849 = 10'h351 == idx ? $signed(-12'sh577) : $signed(_GEN_848); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_850 = 10'h352 == idx ? $signed(-12'sh56f) : $signed(_GEN_849); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_851 = 10'h353 == idx ? $signed(-12'sh567) : $signed(_GEN_850); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_852 = 10'h354 == idx ? $signed(-12'sh55f) : $signed(_GEN_851); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_853 = 10'h355 == idx ? $signed(-12'sh557) : $signed(_GEN_852); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_854 = 10'h356 == idx ? $signed(-12'sh54f) : $signed(_GEN_853); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_855 = 10'h357 == idx ? $signed(-12'sh547) : $signed(_GEN_854); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_856 = 10'h358 == idx ? $signed(-12'sh53f) : $signed(_GEN_855); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_857 = 10'h359 == idx ? $signed(-12'sh537) : $signed(_GEN_856); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_858 = 10'h35a == idx ? $signed(-12'sh52f) : $signed(_GEN_857); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_859 = 10'h35b == idx ? $signed(-12'sh527) : $signed(_GEN_858); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_860 = 10'h35c == idx ? $signed(-12'sh51f) : $signed(_GEN_859); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_861 = 10'h35d == idx ? $signed(-12'sh517) : $signed(_GEN_860); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_862 = 10'h35e == idx ? $signed(-12'sh50f) : $signed(_GEN_861); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_863 = 10'h35f == idx ? $signed(-12'sh507) : $signed(_GEN_862); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_864 = 10'h360 == idx ? $signed(-12'sh4ff) : $signed(_GEN_863); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_865 = 10'h361 == idx ? $signed(-12'sh4f7) : $signed(_GEN_864); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_866 = 10'h362 == idx ? $signed(-12'sh4ef) : $signed(_GEN_865); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_867 = 10'h363 == idx ? $signed(-12'sh4e7) : $signed(_GEN_866); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_868 = 10'h364 == idx ? $signed(-12'sh4df) : $signed(_GEN_867); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_869 = 10'h365 == idx ? $signed(-12'sh4d7) : $signed(_GEN_868); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_870 = 10'h366 == idx ? $signed(-12'sh4cf) : $signed(_GEN_869); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_871 = 10'h367 == idx ? $signed(-12'sh4c7) : $signed(_GEN_870); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_872 = 10'h368 == idx ? $signed(-12'sh4bf) : $signed(_GEN_871); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_873 = 10'h369 == idx ? $signed(-12'sh4b7) : $signed(_GEN_872); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_874 = 10'h36a == idx ? $signed(-12'sh4af) : $signed(_GEN_873); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_875 = 10'h36b == idx ? $signed(-12'sh4a7) : $signed(_GEN_874); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_876 = 10'h36c == idx ? $signed(-12'sh49f) : $signed(_GEN_875); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_877 = 10'h36d == idx ? $signed(-12'sh497) : $signed(_GEN_876); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_878 = 10'h36e == idx ? $signed(-12'sh48f) : $signed(_GEN_877); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_879 = 10'h36f == idx ? $signed(-12'sh487) : $signed(_GEN_878); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_880 = 10'h370 == idx ? $signed(-12'sh47f) : $signed(_GEN_879); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_881 = 10'h371 == idx ? $signed(-12'sh477) : $signed(_GEN_880); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_882 = 10'h372 == idx ? $signed(-12'sh46f) : $signed(_GEN_881); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_883 = 10'h373 == idx ? $signed(-12'sh467) : $signed(_GEN_882); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_884 = 10'h374 == idx ? $signed(-12'sh45f) : $signed(_GEN_883); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_885 = 10'h375 == idx ? $signed(-12'sh457) : $signed(_GEN_884); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_886 = 10'h376 == idx ? $signed(-12'sh44f) : $signed(_GEN_885); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_887 = 10'h377 == idx ? $signed(-12'sh447) : $signed(_GEN_886); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_888 = 10'h378 == idx ? $signed(-12'sh43f) : $signed(_GEN_887); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_889 = 10'h379 == idx ? $signed(-12'sh437) : $signed(_GEN_888); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_890 = 10'h37a == idx ? $signed(-12'sh42f) : $signed(_GEN_889); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_891 = 10'h37b == idx ? $signed(-12'sh427) : $signed(_GEN_890); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_892 = 10'h37c == idx ? $signed(-12'sh41f) : $signed(_GEN_891); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_893 = 10'h37d == idx ? $signed(-12'sh417) : $signed(_GEN_892); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_894 = 10'h37e == idx ? $signed(-12'sh40f) : $signed(_GEN_893); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_895 = 10'h37f == idx ? $signed(-12'sh407) : $signed(_GEN_894); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_896 = 10'h380 == idx ? $signed(-12'sh400) : $signed(_GEN_895); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_897 = 10'h381 == idx ? $signed(-12'sh3f8) : $signed(_GEN_896); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_898 = 10'h382 == idx ? $signed(-12'sh3f0) : $signed(_GEN_897); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_899 = 10'h383 == idx ? $signed(-12'sh3e8) : $signed(_GEN_898); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_900 = 10'h384 == idx ? $signed(-12'sh3e0) : $signed(_GEN_899); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_901 = 10'h385 == idx ? $signed(-12'sh3d8) : $signed(_GEN_900); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_902 = 10'h386 == idx ? $signed(-12'sh3d0) : $signed(_GEN_901); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_903 = 10'h387 == idx ? $signed(-12'sh3c8) : $signed(_GEN_902); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_904 = 10'h388 == idx ? $signed(-12'sh3c0) : $signed(_GEN_903); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_905 = 10'h389 == idx ? $signed(-12'sh3b8) : $signed(_GEN_904); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_906 = 10'h38a == idx ? $signed(-12'sh3b0) : $signed(_GEN_905); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_907 = 10'h38b == idx ? $signed(-12'sh3a8) : $signed(_GEN_906); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_908 = 10'h38c == idx ? $signed(-12'sh3a0) : $signed(_GEN_907); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_909 = 10'h38d == idx ? $signed(-12'sh398) : $signed(_GEN_908); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_910 = 10'h38e == idx ? $signed(-12'sh390) : $signed(_GEN_909); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_911 = 10'h38f == idx ? $signed(-12'sh388) : $signed(_GEN_910); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_912 = 10'h390 == idx ? $signed(-12'sh380) : $signed(_GEN_911); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_913 = 10'h391 == idx ? $signed(-12'sh378) : $signed(_GEN_912); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_914 = 10'h392 == idx ? $signed(-12'sh370) : $signed(_GEN_913); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_915 = 10'h393 == idx ? $signed(-12'sh368) : $signed(_GEN_914); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_916 = 10'h394 == idx ? $signed(-12'sh360) : $signed(_GEN_915); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_917 = 10'h395 == idx ? $signed(-12'sh358) : $signed(_GEN_916); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_918 = 10'h396 == idx ? $signed(-12'sh350) : $signed(_GEN_917); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_919 = 10'h397 == idx ? $signed(-12'sh348) : $signed(_GEN_918); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_920 = 10'h398 == idx ? $signed(-12'sh340) : $signed(_GEN_919); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_921 = 10'h399 == idx ? $signed(-12'sh338) : $signed(_GEN_920); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_922 = 10'h39a == idx ? $signed(-12'sh330) : $signed(_GEN_921); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_923 = 10'h39b == idx ? $signed(-12'sh328) : $signed(_GEN_922); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_924 = 10'h39c == idx ? $signed(-12'sh320) : $signed(_GEN_923); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_925 = 10'h39d == idx ? $signed(-12'sh318) : $signed(_GEN_924); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_926 = 10'h39e == idx ? $signed(-12'sh310) : $signed(_GEN_925); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_927 = 10'h39f == idx ? $signed(-12'sh308) : $signed(_GEN_926); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_928 = 10'h3a0 == idx ? $signed(-12'sh300) : $signed(_GEN_927); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_929 = 10'h3a1 == idx ? $signed(-12'sh2f8) : $signed(_GEN_928); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_930 = 10'h3a2 == idx ? $signed(-12'sh2f0) : $signed(_GEN_929); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_931 = 10'h3a3 == idx ? $signed(-12'sh2e8) : $signed(_GEN_930); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_932 = 10'h3a4 == idx ? $signed(-12'sh2e0) : $signed(_GEN_931); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_933 = 10'h3a5 == idx ? $signed(-12'sh2d8) : $signed(_GEN_932); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_934 = 10'h3a6 == idx ? $signed(-12'sh2d0) : $signed(_GEN_933); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_935 = 10'h3a7 == idx ? $signed(-12'sh2c8) : $signed(_GEN_934); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_936 = 10'h3a8 == idx ? $signed(-12'sh2c0) : $signed(_GEN_935); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_937 = 10'h3a9 == idx ? $signed(-12'sh2b8) : $signed(_GEN_936); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_938 = 10'h3aa == idx ? $signed(-12'sh2b0) : $signed(_GEN_937); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_939 = 10'h3ab == idx ? $signed(-12'sh2a8) : $signed(_GEN_938); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_940 = 10'h3ac == idx ? $signed(-12'sh2a0) : $signed(_GEN_939); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_941 = 10'h3ad == idx ? $signed(-12'sh298) : $signed(_GEN_940); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_942 = 10'h3ae == idx ? $signed(-12'sh290) : $signed(_GEN_941); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_943 = 10'h3af == idx ? $signed(-12'sh288) : $signed(_GEN_942); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_944 = 10'h3b0 == idx ? $signed(-12'sh280) : $signed(_GEN_943); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_945 = 10'h3b1 == idx ? $signed(-12'sh278) : $signed(_GEN_944); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_946 = 10'h3b2 == idx ? $signed(-12'sh270) : $signed(_GEN_945); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_947 = 10'h3b3 == idx ? $signed(-12'sh268) : $signed(_GEN_946); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_948 = 10'h3b4 == idx ? $signed(-12'sh260) : $signed(_GEN_947); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_949 = 10'h3b5 == idx ? $signed(-12'sh258) : $signed(_GEN_948); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_950 = 10'h3b6 == idx ? $signed(-12'sh250) : $signed(_GEN_949); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_951 = 10'h3b7 == idx ? $signed(-12'sh248) : $signed(_GEN_950); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_952 = 10'h3b8 == idx ? $signed(-12'sh240) : $signed(_GEN_951); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_953 = 10'h3b9 == idx ? $signed(-12'sh238) : $signed(_GEN_952); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_954 = 10'h3ba == idx ? $signed(-12'sh230) : $signed(_GEN_953); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_955 = 10'h3bb == idx ? $signed(-12'sh228) : $signed(_GEN_954); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_956 = 10'h3bc == idx ? $signed(-12'sh220) : $signed(_GEN_955); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_957 = 10'h3bd == idx ? $signed(-12'sh218) : $signed(_GEN_956); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_958 = 10'h3be == idx ? $signed(-12'sh210) : $signed(_GEN_957); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_959 = 10'h3bf == idx ? $signed(-12'sh208) : $signed(_GEN_958); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_960 = 10'h3c0 == idx ? $signed(-12'sh200) : $signed(_GEN_959); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_961 = 10'h3c1 == idx ? $signed(-12'sh1f8) : $signed(_GEN_960); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_962 = 10'h3c2 == idx ? $signed(-12'sh1f0) : $signed(_GEN_961); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_963 = 10'h3c3 == idx ? $signed(-12'sh1e8) : $signed(_GEN_962); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_964 = 10'h3c4 == idx ? $signed(-12'sh1e0) : $signed(_GEN_963); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_965 = 10'h3c5 == idx ? $signed(-12'sh1d8) : $signed(_GEN_964); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_966 = 10'h3c6 == idx ? $signed(-12'sh1d0) : $signed(_GEN_965); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_967 = 10'h3c7 == idx ? $signed(-12'sh1c8) : $signed(_GEN_966); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_968 = 10'h3c8 == idx ? $signed(-12'sh1c0) : $signed(_GEN_967); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_969 = 10'h3c9 == idx ? $signed(-12'sh1b8) : $signed(_GEN_968); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_970 = 10'h3ca == idx ? $signed(-12'sh1b0) : $signed(_GEN_969); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_971 = 10'h3cb == idx ? $signed(-12'sh1a8) : $signed(_GEN_970); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_972 = 10'h3cc == idx ? $signed(-12'sh1a0) : $signed(_GEN_971); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_973 = 10'h3cd == idx ? $signed(-12'sh198) : $signed(_GEN_972); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_974 = 10'h3ce == idx ? $signed(-12'sh190) : $signed(_GEN_973); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_975 = 10'h3cf == idx ? $signed(-12'sh188) : $signed(_GEN_974); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_976 = 10'h3d0 == idx ? $signed(-12'sh180) : $signed(_GEN_975); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_977 = 10'h3d1 == idx ? $signed(-12'sh178) : $signed(_GEN_976); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_978 = 10'h3d2 == idx ? $signed(-12'sh170) : $signed(_GEN_977); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_979 = 10'h3d3 == idx ? $signed(-12'sh168) : $signed(_GEN_978); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_980 = 10'h3d4 == idx ? $signed(-12'sh160) : $signed(_GEN_979); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_981 = 10'h3d5 == idx ? $signed(-12'sh158) : $signed(_GEN_980); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_982 = 10'h3d6 == idx ? $signed(-12'sh150) : $signed(_GEN_981); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_983 = 10'h3d7 == idx ? $signed(-12'sh148) : $signed(_GEN_982); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_984 = 10'h3d8 == idx ? $signed(-12'sh140) : $signed(_GEN_983); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_985 = 10'h3d9 == idx ? $signed(-12'sh138) : $signed(_GEN_984); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_986 = 10'h3da == idx ? $signed(-12'sh130) : $signed(_GEN_985); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_987 = 10'h3db == idx ? $signed(-12'sh128) : $signed(_GEN_986); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_988 = 10'h3dc == idx ? $signed(-12'sh120) : $signed(_GEN_987); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_989 = 10'h3dd == idx ? $signed(-12'sh118) : $signed(_GEN_988); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_990 = 10'h3de == idx ? $signed(-12'sh110) : $signed(_GEN_989); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_991 = 10'h3df == idx ? $signed(-12'sh108) : $signed(_GEN_990); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_992 = 10'h3e0 == idx ? $signed(-12'sh100) : $signed(_GEN_991); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_993 = 10'h3e1 == idx ? $signed(-12'shf8) : $signed(_GEN_992); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_994 = 10'h3e2 == idx ? $signed(-12'shf0) : $signed(_GEN_993); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_995 = 10'h3e3 == idx ? $signed(-12'she8) : $signed(_GEN_994); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_996 = 10'h3e4 == idx ? $signed(-12'she0) : $signed(_GEN_995); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_997 = 10'h3e5 == idx ? $signed(-12'shd8) : $signed(_GEN_996); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_998 = 10'h3e6 == idx ? $signed(-12'shd0) : $signed(_GEN_997); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_999 = 10'h3e7 == idx ? $signed(-12'shc8) : $signed(_GEN_998); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1000 = 10'h3e8 == idx ? $signed(-12'shc0) : $signed(_GEN_999); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1001 = 10'h3e9 == idx ? $signed(-12'shb8) : $signed(_GEN_1000); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1002 = 10'h3ea == idx ? $signed(-12'shb0) : $signed(_GEN_1001); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1003 = 10'h3eb == idx ? $signed(-12'sha8) : $signed(_GEN_1002); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1004 = 10'h3ec == idx ? $signed(-12'sha0) : $signed(_GEN_1003); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1005 = 10'h3ed == idx ? $signed(-12'sh98) : $signed(_GEN_1004); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1006 = 10'h3ee == idx ? $signed(-12'sh90) : $signed(_GEN_1005); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1007 = 10'h3ef == idx ? $signed(-12'sh88) : $signed(_GEN_1006); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1008 = 10'h3f0 == idx ? $signed(-12'sh80) : $signed(_GEN_1007); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1009 = 10'h3f1 == idx ? $signed(-12'sh78) : $signed(_GEN_1008); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1010 = 10'h3f2 == idx ? $signed(-12'sh70) : $signed(_GEN_1009); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1011 = 10'h3f3 == idx ? $signed(-12'sh68) : $signed(_GEN_1010); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1012 = 10'h3f4 == idx ? $signed(-12'sh60) : $signed(_GEN_1011); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1013 = 10'h3f5 == idx ? $signed(-12'sh58) : $signed(_GEN_1012); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1014 = 10'h3f6 == idx ? $signed(-12'sh50) : $signed(_GEN_1013); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1015 = 10'h3f7 == idx ? $signed(-12'sh48) : $signed(_GEN_1014); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1016 = 10'h3f8 == idx ? $signed(-12'sh40) : $signed(_GEN_1015); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1017 = 10'h3f9 == idx ? $signed(-12'sh38) : $signed(_GEN_1016); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1018 = 10'h3fa == idx ? $signed(-12'sh30) : $signed(_GEN_1017); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1019 = 10'h3fb == idx ? $signed(-12'sh28) : $signed(_GEN_1018); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1020 = 10'h3fc == idx ? $signed(-12'sh20) : $signed(_GEN_1019); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1021 = 10'h3fd == idx ? $signed(-12'sh18) : $signed(_GEN_1020); // @[direct_digital_synthesizer.scala 67:{8,8}]
  wire [11:0] _GEN_1022 = 10'h3fe == idx ? $signed(-12'sh10) : $signed(_GEN_1021); // @[direct_digital_synthesizer.scala 67:{8,8}]
  assign io_B = 10'h3ff == idx ? $signed(-12'sh8) : $signed(_GEN_1022); // @[direct_digital_synthesizer.scala 67:{8,8}]
  always @(posedge clock) begin
    if (reset) begin // @[direct_digital_synthesizer.scala 35:22]
      phase <= 32'h0; // @[direct_digital_synthesizer.scala 35:22]
    end else begin
      phase <= _phase_T_1; // @[direct_digital_synthesizer.scala 39:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  phase = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
