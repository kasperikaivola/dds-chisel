../chisel/verilog/direct_digital_synthesizer.v